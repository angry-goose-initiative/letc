/*
 * File:    letc_top.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module letc_top
    import letc_pkg::*;
(
    input   logic   clk,
    input   logic   rst_n

    //TODO other ports

);

core_top core_top_instance (.*);

//TODO all of the inner goodness

endmodule : letc_top
