../../rtl/letc/letc_pkg.svh