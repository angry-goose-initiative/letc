../../../smoke_tb.sv