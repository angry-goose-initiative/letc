/**
 * File    smoke_tb.sv
 * Brief   Empty testbench for smoketests
 * 
 * Copyright:
 *  Copyright (C) 2024 John Jekel
 * See the LICENSE file at the root of the project for licensing info.
 *
*/

/* ------------------------------------------------------------------------------------------------
 * Module Definition
 * --------------------------------------------------------------------------------------------- */

module smoke_tb;

//Just end the simulation immediately
initial begin
    $finish;
end

endmodule : smoke_tb
