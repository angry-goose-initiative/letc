/*
 * File:    letc_pkg.svh
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

package letc_pkg;

    /*package mem_pkg;
    //TODO perhaps move this to a different file?
    endpackage
    */


    //TODO

endpackage : letc_pkg
