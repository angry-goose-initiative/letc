/**
 * File    learning_tb.sv
 * Brief   Testbench for learning (System)Verilog!
 * 
 * Copyright:
 *  Copyright (C) 2024 Juan Segovia
 *  Copyright (C) 2024 John Jekel
 * See the LICENSE file at the root of the project for licensing info.
 *
*/

/* ------------------------------------------------------------------------------------------------
 * Module Definition
 * --------------------------------------------------------------------------------------------- */

//TODO the rest
