//TODO like amd_bram but width must be multiple of 8 and we support write byte enables
