//TODO add structs for between the various stages
