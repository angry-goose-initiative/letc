/*
 * File:    core_gen_imm.sv
 * Brief:   Generates the immediate value
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module core_gen_imm (
    input clk,
    input rst_n,
    input logic [31:0] instruction,
    output logic [31:0] immediate
    // TODO other ports
);

endmodule : core_gen_imm
