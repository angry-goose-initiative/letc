/* letc.sv
 * By: John Jekel
 *
 * Top module of the LETC SOC
 *
*/

module letc(
    input logic clk,
    input logic rst,

    //TODO what ports will be exposed?

);

//TODO

endmodule
