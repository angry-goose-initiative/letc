/*
 * File:    core_master_control.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module core_master_control
    import letc_pkg::*;
    import core_pkg::*;
(
    input   logic   branch_en,
    output  logic   invalidate_fetch
    //TODO ports
);

//TODO

endmodule : core_master_control
