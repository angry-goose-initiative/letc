/*
 * File:    core_top.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/


module core_top
    import letc_pkg::*;
(
    input clk,
    input rst_n

    //TODO other ports

);

/* ------------------------------------------------------------------------------------------------
 * Connections
 * --------------------------------------------------------------------------------------------- */
reg_index_t rd_index;
word_t rd;
logic rd_write_enable;
reg_index_t rs1_index;
word_t rs1;
reg_index_t rs2_index;
word_t rs2;

/* ------------------------------------------------------------------------------------------------
 * Module Instantiations
 * --------------------------------------------------------------------------------------------- */
core_control  core_control_instance (.*);
core_alu      core_alu_instance     (/*TODO*/);
core_gen_imm  core_gen_imm_instance (/*TODO*/);
core_reg_file core_reg_file_instance(.*);
core_mmu      core_mmu_instance     (/*TODO*/);

endmodule : core_top
