/*
 * File:    core_s2_comparator.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module core_s2_comparator
    import letc_pkg::*;
    import core_pkg::*;
(
    input   cmp_op_e    cmp_operation,
    input   word_t      rs1_ff,
    input   word_t      rs2_ff,
    output  logic       branch_en
);

//TODO

endmodule : core_s2_comparator
