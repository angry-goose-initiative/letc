../../rtl/letc/core/core_pkg.svh