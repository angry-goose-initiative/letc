/*
 * File:    coraz7_top.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module coraz7_top
    //import letc_pkg::*;
(
    //TODO ports
);

/* ------------------------------------------------------------------------------------------------
 * Connections
 * --------------------------------------------------------------------------------------------- */

input   logic   clk;
input   logic   rst_n;

/* ------------------------------------------------------------------------------------------------
 * Module Instantiations
 * --------------------------------------------------------------------------------------------- */

letc_top letc_top_inst (.*);

endmodule : coraz7_top
