../../smoke_tb.sv