../../rtl/letc/limp_pkg.svh