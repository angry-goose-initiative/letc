/*
 * File:    TODO.sv
 * Brief:   TODO
 *
 * Copyright:
 *  Copyright (C) TODO-TODO TODO
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

/* ------------------------------------------------------------------------------------------------
 * Subdivision
 * --------------------------------------------------------------------------------------------- */
