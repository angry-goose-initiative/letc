/*
 * File:    core_s1_control.sv
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

module core_s1_control
    import core_pkg::*;
(
    input clk,
    input rst_n

    //TODO other ports

);


endmodule : core_s1_control
