/*
 * File:    letc_pkg.svh
 * Brief:   TODO
 *
 * Copyright (C) 2023 John Jekel and Nick Chan
 * See the LICENSE file at the root of the project for licensing info.
 *
 * TODO longer description
 *
*/

package letc_pkg;

typedef logic [33:0] paddr_t;
typedef logic [31:0] word_t;
typedef logic [15:0] halfword_t;
typedef logic [7:0]  byte_t;

endpackage : letc_pkg
