//TODO just instanciate an SRAM module within.
